module abs(In, Out); // 