`define GOT_UPE_POPSIGNV
module abs(In, Out); // 

endmodule